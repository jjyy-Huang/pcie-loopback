`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
T0IMb0CNHGINngqK01lEyA7aS9ZxSWrBhNV1CS75TK+6mjV9T9Bsvp2+Y23w7o3ZhyzJUa54DYER
LaRX1+k3iT73pW4AZ8gWDncBuT+1L9EwgBZekiwwqaiwRAFy01+/6eNNMR1V0ebF/0EUX/bSxk1N
GDi2QR04mEHUO8XG/qf9F+G5Of4b+xzXnYLLSsrsEWbEyQLKOmRvq8Tfh6ziI3Bx42fXvVuEuv22
w0b3VYNz9ggsVf+yFKYjNhfOgQW/FkFb6FdDb/2atESkWzfT7xnH8tylAwttYGJ+qjDeaK1VBqBJ
2zQOUO9h/Pggonze4YVeq/bRLQZvuPJOiZ/mrw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
xrp5LA+VLb5YVvNodgQE83sioHSAEy/UaW9TZMPkpxcK3ERIlmirtYO2Ju3owSK1MoT7XrttYdzp
7hCHw/UPjR/5HVii8Zk7wwyaEgjzgekskXVPmqo1MQg83IkgDa13CLQhA4m0Sd4Ly2twiInvzE5z
r7DPh0CE/v3B60xfGTWTQhchtozW2okSt/fkqf4hJg3UQgPFcXIJTTIAZcn5t9Ank+uFjHM5dz6Q
vxtVxH/NVF/tcCiiZsfxTkWfrqjrQLB8I2+kc010n3NvWB7hffX0HaVzL7ehcJMI50t7eOogsQG3
KCcrhmFSa0CjquTzBnmeA0o7iX/FaxCcb5KZ9gAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
IVxTgbfCcOtLBUZxStz4VBabWnBUXTsPT9pBgI4pGUjDLj5NHu8oM3FygJbp+eFjghj3Y5CwYYyC
sZ1ZqXQaEw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
byjpmFziiyeqVYJu1rGpl1gCdm5YONbq56+GoFfsBrPEBzw75Bp6TmQadOuRQv3AjiDB8NvqS0G6
nXiI8ErVX1Bye3Ra6V/ytQsM9D+ccJMp8603LkD2Aq2cc2EJ+yx5YH9oqgv5yvUJ4u197fn/7fao
xtZj5zJUfthoYX5nsJshEOiX7/xyLHyvI2cD+2gjhlo8gEqtuYN9+Vto4eUEA65mex/GxdFFwfDS
/zrIbKtQxBWjq+hqSL04qgHiGqQPHJVzQV9G/h6eFaSijbmnweeh2dTOWTn44qolgx43KHNP7GJ9
woccnUzpRcJPBw6lHyGN7ziRuY2N2S6kJWIsCQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YSWGWXuE/aeckYnoMYl+mumdOZE7vWAxciFOegsvpBU6DQXt+gpNNxVf/IJ/ICCRzt6iZ9epMFnb
xirQC/I6ChRtvZoQoCTH9WQbqdmMB0yxZiLIHSZ0sUJikQOTDUOJAaer6gNFGc/cHWBhXGokhHwy
fkDVANFyQ6Z61Tu+IhoInyAaXqDzCpwTUKZuf+xibxd9YBkVzgNxs+GmjuPR+Ew+YqXv4We4Y+ex
Yi6bDjYSe33bnr30UJuxykOR6FcCkfoAxOcpQ2dQxB4tSnc1UmMywjHjDhVW+yq9vEQk9CV3LxBN
I81MpbrkX035HeahNpHTDupj+iIn0Kxs6j9eRw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fB6nSZGZqlep0wyeW+bu9jq0uEHtpEDXVq4ezvVlhHaRZYd++gOSljRM01XdnueZWb5AEHdXFh9a
Hyw+UWNhMx+Lu8cVO2ZoE6F+G2xrTbFDQ5T2JNAjZUyKI8+268j4HMTtfpBS2J9u6gKdMCz2Y2hU
hioncjt1iAjYIgz38rE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SCEM2eZgcqBVBNeP6oT6xj6wPa+MBLvNUXg9P4SaHfFoSY9F76sysQe3Za18kyLcW4+p0eHWb8En
uW8K5u2ZFz21s+YDXO0NUJ7SePUq4MSoI9Gvu0lsFVxlEvzH0hT8LdqtyjafIRui4ghwGcARrUMv
TgXyfU9A35x1QF4z1SLhT73zAvWCwK3Xxm2T2ulrPqx8fBVvBV0BROkNZ14sJD09cwTn7FHClwRy
WHLvgvdMs0a/XugBDbiGTJeBvFG5+e8fD56893d/hjHuuhID+64YYtveUoxBPqi/FUw+WoenYZUB
Kyn0xq5106FkWWT/iGTrbfKOUIwn9YZ43PkX+w==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YcQwcMllQXztRjmMR1478WJve27gD1+sADFNftBucp0KuZiLe+fudYOUWF/2qwp2Y6yLPv7z9OA2
Rn1qkr5XZcQVZOOA7aajl4v6rAlYaQMZk7XtaeF8uu+OOkd9KYD8tLXq/QjPVPhqRyJn4peHqPcw
9ltGFB+ILXtnqY1Bw8YFHd7sSw5jSiUThG9bfr8CG0UERwhw3tr8kEHYulWQschLO2Ug5FSPD8ln
zNKtbDkpZxhBvYiHwCypaEXOSwJjpGr9YeMgnrArUgyZHjyRsSOEBQ/XdSCz+UoA+OSL4EX9Out4
Lyjr0RmHxBXn80loxTvAZR5Iew4o3DndiOnOqw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AXS+RAjxe+pQllXoc48TQm2q4uLBQuu1Rzn2tztPJPReQPAKTSKbTYDeFdDRlp2dgks/mtMjy7Yi
15A++LkCpvCNk5EBHRbGfP5Vh2dBoJ1TlzS0I94XuT9rgx8VZLXivYsSr/Q+lSLwMT3CG4OVnjXO
GoOo7VDkhvSbD7kdsM8=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N+5zSkl/Uzt/qSVmd9UvnkyO1bO59o+A95aZEJWoetkt9q0yPl4iwIJPrEpfRxncUVYT6nzc4TCT
+npKGFCil49RK/2AKGV6odNs+DyWrJ6u/JNlfdjkJXajxYNnnYA0rD815lt35kVrYy30NVRR04W0
iUdY/CTBPxwJMKzuHNkOvP85NDXL4sXT2EIK0z/bofjzDQCTGaUs3Km0brlOxXLe5isuI28gutTo
bF+gvnRNagY3Drg4bpWEq+miS/CBj+9YuOs3FjEqwDb2kPHYU9l7bp4sDkxMePiQ4h4tGVMgLT6X
4e0HR2dQnW6X/6RWpas8SVrFmbnFT42FiNDDoQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
Sj0OUBcYhR8Nt3DxgVDF6uYYhfqOFrcDEgEDaJuLsMvlvhaObSJ4Kh0jQc73iz+2/3EXlk3MEKQ1
kxiaN6zh9jqaZlPea4/48U5qjSoJ9SF/ZgVPGf1ClVIyAw59UoKJeG9mDN8PrdeD/jvXl4l68kuD
LTZ33sjHr4r/+LotGE3WJbCorCXfVJGHKuzFhRjLdRl7IGqSNgahvJdwZYMwihC3xrzJAZZW4dkE
EoHOjbXL92WaRKj/3qisJ6fBDslsRxaBG5KWEScOXw6y2em8H6u0WiFPpJM+rFa2pWp2NMPDM2nl
9v85n2zD9mR5L0i6wF/NqSkZWI/x2kpZFX6UGuj2c3srU3B6vdHnsqnNlc3cZ/EvyMFhIYHUaKpe
UZBvQRZWhnvd1Tyadr4dcO+s1tlPnSX0pTkIkVu0CrdvfSIO2qrNAxX7coRincPgQylNJktoekSX
ClRsy3UKM4AKj+Q+JaJAoMSteBYyWcYUxO4lFNb34oVKsqsaiRp+4YFV8qcdSG/0db2KA1XCLNzh
nahGA+nWtwQmaSnbdCmY/7kVbrw39HwKyqLQ13j2z/IQ3dIR+pVZ8EY4LuyUbzeTKh9LnV2oKup6
IvZ3HZFu2KJpPp9kYH9CzrWDyZAOSHjb/gwqdyM+ixrKyXAC8r1usenkCeIzjO6Zn/cXbfN9wQXU
dDI11YRHJmWrmq3gqLJg0cjLI4RcDIhMmj9FFdrAMYoS8JctEh/stplg6G1CjhzVvoer+xHY6LUD
K9bwhezxAJSMXPPVNu1S5N7hew5/vKTVnjJoxwsiFkx7MRAAsfO3eM9U+xbpDLCnpBzQUh1Su4/K
rWCV8mWFgSDcVOemL/7MXGt1Mv8qcLgOGxUxbTgq5vQX0ygr5JKh+nDXMpjclt/qAu+eiQ10MIUG
X47tXqVpzTnVY0YZvIxACrtUuzbsLG1k41V9OJJnVYKSVcZ8v+d9TJaOlsnhYulga4JbpPCD9h0E
uYqFQaSNrwhiQZq4f5jOy+bQTLJXZ2hziJ4Wj4goG5woHOzbmOY1hsNf+M0BgACD91LgXN3391od
8YqOthkbkLY5USQtJWYz7tmw6OFiZ0SZncLtKfejK+MdauelxFLLAPNQqDB50KC81HXobdOAK0O8
pF9Y4YtMXFtqaWR0H2IxKj6bp3V6yHIq2a0hBUKDLJg5L7vnGN8YIlD6aHt1vDkAYksk/DTFDFh3
yrHMrUJrAP2e7r6FalMG0+rYXHeoxfhZC+Yk/MlLZw/HRcIohwFW6DK949sWp9sy2R62QDdJ29qF
1ASH1rWwWu7siyJ1rsO9pYBEh8rQD7snbUfTOB8TDJASWm64Fh8ng8Q+K0lnrnhoq8Yf0IFqwTC1
tjfFWrspHyyhOks43OipxhP0EYWvIpDJijfzB69iLuV/dbZvy0fKJi84VHwDVTBSgWrJhKNT8ak5
tU3Tb+7dqyab/68mg0qDnTo0M0V25/vJBtI4yrYpqAR+CqDSHAnD1sMjWLcSdzabrjeRADZd/BWK
+Jq0ZruYA8dae7xMlTqzG6bSbPx83UMljc4Nl1Cp84dEmzNniSfjhrcWaj8ikTcgKWZReFZELSUu
N4na9yeSPkwwMsLMs4iItYhX3N8QkF1lWX7mPTprJidudRn/sm7c8r5C86wqEvzw5Y/YWnZKtgto
s4AQa+BmSmIcMk5q5dXP4UoplCNSGJ29Wam43MZXt7zps0jV2CK6cq12WEVx+arHNSHhPJTOVA6M
oA+nFgd/fT++1Cq6KwmrzlT/HUd8ce7v0RUiOv+mwkV9QW16FbTkvcji47ZzOwemLo1IBg7uOnZJ
NZ35xKOlQpXxH45M3e/bT0Cd1ANxYQhKMwc47acEDw2G6QMXe61ERk3VIiznqSDBs6WoXTsp41OY
vK6mi8QwgoDB4C9IO2pUbZooQN3uTUB4Una0ocrNnpOaZPRhvHUetm6yor8H1onfwyxjlMtEuuXr
3E+TfQNDg09wMrmnMxs932OBUcxm5qpUexA8yi4gvRgIAxJLGv3rhvOTeUyyj0g9dIUwlLuVq/7h
vOLja1QF61QKJfl8vFDBWG3YITObsttpAVScjYZqIE4nwLUyxY2yT0GLmwC+/NYTZEj0kvy1+lTC
WeSVR6tVkT25ov++nqv67JIDK/WCTfkfOohXVa4qJdIfL0geSHNdTEAJG8YNpntPlkA4rfOR6TBW
jEskhWbWzVhyqA1zZA/Kb7BN6m/BuHKfBg6ZFPWFllDvFYjcL78GKHO2OyzWiSMZ2tBaMMxtYfqC
UfLj6rTSQYie7MHUWRSTfPnB1NzdhBtIOhd8Yt4WTiQaw92qYxczt4onxppmef6TIkh/bVDso1mI
oe1xNDZjHK9vz09JyKyOg18DI4LuU7gen3vF/f+SpfnL7ewSEoLQr/Hl/Gh2ZugS+ETm/p4jv8vD
BQfqDn6GrW6eXSzcUKfo74cvzKIo+j5pgQ56OZh8qd1BUJ8a5apzgmR+la/t/xqMybjFN5IIRNAF
3sDQwaNNZBWZDi3MfgzaeUJvW9xsdrMIClxKaXipmiSlNn8S6TJtFvEdo6CMo8orE3hmg4aXcYFu
Vl1PBh7Wg4hUREpUF6KFEw9gIaw7Y2weK5KL8Wbh4J0b+MV0d+egN1UUo5DSe5xTucn3/VYU1eD5
tCGj/8Dz43cSHtFmyItayIX9MN1MP3ROha9hmGJycIV4dlyKYquRbfAYhEjJzwjkxNQVNIKHbgIY
3HcN5Y+uwW/v801DDyXHapDl4Yi9axrxNikgUdzynG+yKyThhZuyQu7eQCin+LRP6dxLYBi7joLt
PF2rnw43HhbIDSQtC22sIvNKva2vV3Pi/c7XVDfpyb4lc9+OKZBzg0mEOmJ2cKDbU22KnSRc921z
bFHUZ3fjDmBq7H+JMv74ELH0SyhGR92b27gsKarFQ3ew9XN2/YUsW6wlMljYMeBAQzJ2RAKwum8+
o7TsgknAeqDmakslXWqEmymlioyaj8MohVkfFwY6hoAHgc0KXkdXTPwTN0QRy3nnjSsePt4h6nAW
O+FUlr5JLzylDEM4pgxMDjvixv+ljkvCoAYwkryVJtHkjzfPbzFUUAGjkhEH9uCdTNxUaf0QJIfc
uFDbV08CY8xCAxBHqEGPDE5CSNGoSxllnlvjN8+58NqZ59qdmicX71dxk4quljs5ShXLyBUfFqq6
6/viF8zcYZK630SNM/HVm8P/Ifl+Kk7DuVHmmHTpeFoCIuLomT45kYjvi78Dz/LIFyXBjiH8a04N
biZO/d0dCN3ztN2vaNAsoXoJmrKW1319RJ1S0rbpf8x/B8VzGbuFaW1T8mfmgJqDHHdP9tbaJKzK
xmdQ5H+U0lYElRVfXu6wu3oyyCvKtytARCkxux/r5jUCVetWIAXxbNarmT0CJ0CcxXrbRgIGtLUZ
YCPoLstg9nJ5xC7kbCGfnGsoR92CPOffLeJmyOV4+Hjz6Ux9jtNRARa9mdWtxwvaGpcY69F8sUwT
ChkOw2Kv2iyZxpoG7xg7nd21AEooLIC81KxFMZqY2UGs4kL9LYXbef06kVBXL1yqVETosol2ic2x
ds3YcAlqRNRfXdvfbeZEm2BkkpDEa64J25ogAXKMaewecP1dT2Nva7VZfSHA535uYqFRruSLAgAZ
3YJ5BVplnb1K4FJowCydaoZVQK+3zTGpB22S7Li3VMgHYPyYCJ02ujmDXHPuMayJo0ywt4onKaKX
HEJpFI1L/B1UUUIMRTDLHwdJ+tz5DYoe69iAaQT/rkbIFiziGrcTSNSN2sPO1qUN0CkPd3ms5ftz
5xyFyn/74Tq3ba9GN637hvCTZVEEgN2PIWsOwCTWcZ1cb0l/Ll9VzIwVkjiBJVDWAtuog30aDq6p
E7CWUBkj/NCwQQFn06nGDDmcs7eM64nremVEqEWqT+ZifonHqQJ2L0/YF+2sGjVzhIj+N4TUkAZ6
iYvkvCVRoypqSwg6HCtHRDZz3tWvdrPcS9qQgu+zl9+ID6Nd4WpxINwZSF/j2NVf5MJCY1C64tM5
j9TX8a6FiT0zFT3+Ygn3psn9dQgI0XKOnKvoNXwvfyDJgvuSaff7AVCt1GXfOSyOtFgOANZivipd
sqHemzl9uVSHfvQ/QDuoGthSYPKCzOgtenZA+xFxZAMNGHRaTn6TiTMINJ3gyHHTp75Pa9vq4Iy3
XqVT87KDsQK1fU3YSyPNbhUy87Ydu6XnuvdqKjarodAERQI7enG//a8QE8hpyrhbgi+lMPGNwWrv
niKI96spFRK9TllkVdhpCfbXXVYX8UAn35ixZJYAaIe8zdXYAHtljj6HLfvCh76zFO1RBXN1jPno
VPmgjjUsAENqWkIxrwf6bW77cucweqzagArbI0ZlS0w1/FwgMrvsiFSDKNSyUyy+5kHYYjF3D52y
k7owWew6rCQNPSO8S7iaFDkWtclarG6Z38RC2f32ef+neavbASOJjt4nOk4j87O6fmKkobRFK/+M
xIy2pWlWZZH/Ntz7yg9YTL7k6MDTMODxGAau5+wlqe3Dq3OKigDayEyjRgrK1BuZbnQb62VVmi2g
kMc+zXnUGuO5Ep9jf2MCJg0Rtq3PuKmeRuD5LE5KhS+ruf8XnFVXhMighfszDHxtrPHZMn25EOzT
3cq6qX37HCOlfgANjYbK8r/o2zOltQwdIhBILa24vITxeD66bPdE8mpHAfEKuyIT8chT4YHh4SX4
u6c5khkIDeo9tWEcsogKp+GdFWA5DiZUNo1n//9/DpIWnY8wYP6d28W0SaFp7T4BgWUWE3wW+Ea3
LWxM0OKoCqWfOoDY3puVrtiMEEXJtFdWPBaOfS94uOsBLTjdKBwp1bDgs1bSoMxJjasi9N+1/wxx
0ESVu5fuKDnc2NKYQ4WlNjqD0/eVGngwg3H1X/UFKugThNB1YZqYmcv10OO0GCGrp/xyVegfhOqp
OVDR4U6inUTGP0fpa6W6j0NKj/tavWTGEBCRFv3BhzTJBQokiZPfx5paUtnSMBEKulkXsjIH0ni0
q5IyIPW+/bUYyYEE4l+ZPOLbAAt36g+n38PKGneSqTk53LjEiOHKSMI1xuFKj4yrZFDXIn7woeeE
RoBZoZPTn5vZhlDaGcNiIhYpg6TWnOZFNqybtNbb6PtbqSoUCH3A/mUgCXdR+4hUfvX0CHIaFIh3
4a+uX2/T9J0aZQ03l9FhXhM5hA8sC0oKTMvH0ntejKf3VhyBQQEm5XEjOxoi2vdcMd6RLfDTCB7T
GtlvequIeiwgoXbKcInwmaivlij19DwlFQoC2UrDsOXJ6zd9F+9VomxEgiWG0TTAO9T8Pz5klSv0
G4yQhs3sib+/aRTB7IpmkmZTiJWUe5gzoNdOxv5RWIFNmZAsFv++5jSSGpyFiB7Yvlj0AVNBUHS5
LDmFCtqUBxJOBvJiQiMBe5q414mxUQqAS+tQCvJdASEQtw9aaeIkZADmjpZXm3N0A/AB731pGcNv
vUvSt5H8mkLetpbKCLyRO16Nvyzjgicq/J20myoTpH2aztQJhoWcaEuXI4BpjlTYgIQBs2E6YczT
klx0EWQvjk1bRnXG50qLMCzD7S0Dn0SizI2C5YxhbfmaodMZHKTjeyZwN0oARJvxrRsiITqudoay
PBF1YEgWEjKu1UWcMLS+xMJUd+VPS0pSHKmaRzMTHPpP5RrV3v0rO5u7GishQ+ippdLEjmv6g4pP
ysG3iQBhKU+s5VRFxhnHz9FiAdRQl3opd3cdT5OSS6kQ8ZTI5crlsZV+mg0Ll6hyi2H93fsYUBrA
eEgIw3P/KOigdGWM6AkhAkDOC9B70df6DhSvuIj81aTgDP5LBWgUBcJNmx8DPLPAOLS7bwa+602Y
GaNbrdApRCJCPi+tBLUkZpIx0GfDYNu3ttLxIeDbuplNu6pbaa9hPQcVICYMkut4VCAz14CKN/mD
HfqiFXPEJr19qTSoKmhRuqHyeT2B4Jz5NS935Q0By+yECPsauWlu86+Hk329Rm/X/Uy8RksXdHmN
3wlo8h2LdSueoKBT5uNEGsZQyOInyT4ln1SzXIMQRr1si1ZGKAlAwRs9yUFM2zGN4u/3WV5g4n/r
k2vyIeVLKbU0ewl9ubq9G7CdXgAVGOH0iDsJ49SgzYyDDKckQutVyUMte2jxsjkU54Gs3lDQJfeo
iMGE0X/OWIg8Tbv+X5ziRfwBEDYZms8BVymTO3lM4bpO/QxHNrcvMjnWUgJe5btrpyccMPAQQBoW
ocMajkc2Y/CgJpTS/+kbUg7bL/NWJyINfTgGbjQe4+WUQ8HZ7WFoXAQifRuNDJKwp/DIf7bnc143
dRWwzhhcnoEKm4LmPUk6HNUlGX1n90iz14erZWTDWwGT0u0emottyndd2iulJ4zIAkrN1ejg2s2I
crgzSZm3lWMuSNRRVwY1z2X4qiWAg7iPkFsqepCbjhdIAwULFq2KTTwj8FaBeFiAmLMIHu2b9CGk
W/sWJzry0tEnftge4x7yiAsSiH8cf3a9C7DU/tvBvdUE1r50CpK4gI5LJWrGVQZds68kiCyF1AwZ
73MtmPqMGMN+eG8WkSt3yj3go4zLplaOew/B5KpUDiSc8UyjBPEHrZhOBWDzE7Z30GqxMmw6lo/s
Xdj5LgVyd/O03KzveiMXyJaQVRIf1dbv7XWNs59lYuuhNIdTwutfXL3wf87VbXZBwy70EpHO0bKi
eodBjdJwvBGApsn5F0//jS3ueIFYwZUXAgTQQgqGFWqq72XQIzuoUJG2O/7rGb9hjykOIOpv8cp4
0fJPinRGzBKeJolPVwnZlJR2Ofd5uESSbB7ZiStHUS2E+J2vHKEizSg4ubN7EZmrv41b2Ur6gSH3
0V3P5XcVogoqLvnBMrNaUP4Reg4rNjtN7MI2NRsry4BAx7xTaFqiL1W0LRwXFd3/j7432ag5sgEQ
lb0XIUWE1W/xdn/OiuWaQIvIwI2U0knGWCOoad+6REruPY0+VUYO5SlciKQc7PO3aniooT0Kq1Ge
Foz0ViDbj+3Zk/22iXH8Jgb5FLi8foNCk9TwAnJUn4JkxZHjNgZ9FgHuGl/rp30okWOajCAHqAkE
ay+TYm1KgVUCH8lQGAPd3wzyJEAYMTUXDdCVJ4hS7TLZB2gymCBdouqMLSZWy/R9tr9sKJDqI5qw
7C427U7Oe1gWNQeFq5askStbg0c16QpytT11LYt4h98y6o2fh9sJOAe6wO6TYnLynFmA7DAe4B8G
iNeDcj4nbPrP8bN/0jKwiAqA8F9ekoTcA7TWs3nXspZ7zWwK+KHeKAtmc8yJErpnBi9VOINiG20G
oBumAS2cgZV5FhGVqp6s8RZAewS2XN4V359gM4j+/AIimmLX8vwLys7NqrIDjKrzIBTd+RceH3JH
+M4kSON8ztYGW2q6Dok+85X6QOytXE8fHSHCVaQTCP1XSD4pPIX4/Shgn8mj1wdN7R/y0J/a1/Az
7KKVGenUpg4ja4RqHrpgNWQ//ieHs+vuYIq07qgWEJLiWtbF589+RaOzU3aGwDo1rjPbmcmDcz4/
T9mPn6a9C0EOnCLnAF+emnAw4w8K1JLv1rewllO/Pk11AR/GPz8hhcP0BtZlAIXyeEf8oPPtp/C6
7o4lUGTs8wg5q+ZdVJghHQIVzFX+6B22PPjJ8wx+YF9bmmXDGdWz0yGde7iR1MURNVesGSYToq8w
8ixEoWz3YUZ/GCrFfA+SQZwhdbMfVP089XrTp9WvoOzlG4zh1MS5sn1VESudDbvtORZNhY0uaqVE
4YYIzR/P5PgiNRU+VRg6u6IqkEtshPvfoOMPAsbZKwA26FXJfbxN78WLASjNv69Rkj1pIBc8jyoT
516ESFHu6/H6jThLsYUecInLaZwE+MVTom2v93cDIHG+7/DdSfhZYioFaP5HAUYOI2HVrSPfgaPF
tDJs2xpti+Bv4quwkE2fnxcfJUo5uiI/XUAoXRVeS+/k+gRizbcA1e8BRo1+1hCX/cN/lc40MQ3o
9Aw040lGvz2r9ByA/Xj9rrc5p/AI3eglg9Pc4q+wMtvHqwpL1ztogTzJW5eN2eRgvNTGlLdcCgT4
+RbLN/yvWwicPidoWXsecW0soNSpuk5h+89BCBxenACe4U85W6dCLeMZsavoPX3luBEkPtgryVrK
6Gni9Aj7R02Ls8zJNA8iz1CxJsPZ8/2dDPDjEVddXIb0JZrW6RweoUeDGQR7LL5yK0bJd2e3kq7Y
S9yPqQA8UDJMgH0O4cOKFoE2PbGN6vYhbmlPDBJoIaVly1RskH+pOoreYDkWL02fRo9/W25mQUCE
y1tgAxpy5h0h+14tJpzkCzsfT2QUUqz0/BEDhofhDX8KuJaUelBTNwvycgIKRlH/ETydSRn7vO6Y
B7v5oT5TT24es6cwyj6MVzGL5eePAzxz8TC4tbeJDfpesCBFqrar+9KDWE5Q/uGVNclEKhmiV2pJ
50z3Njas05I4L/RLxK2+dNlUxT11O1ikbDEC4gKJtykuTovJ7ESQLs2hOE2COGU8DiP4XQ1EBOsA
lE9NceFX/N/QqafRTO8aOsdMvswKAgI3iu6UxfTpi6SdYW5MTs3FErGE9ePlNdM5EXuDP4Eva0RH
wGo/jtfLeagQa8d10Q697c7rO7OtuOJ9RDksxVfMlybp8qqtpCsfJr1Y40K19+/phhKMxeNpznO8
FDan57dXsUFKxu+6tz9hg5YfBzuu8UZGonOe4goZo0nIbR/kXtxau5vlvRci+L8WTWdoE+xlip5x
op9Ue6trQeYq90KYw9D+OX+MtS9pkpAFSQMvp+8RjRiKlObse+k0/zqbPfkt7UTTTIJ1DB157f3+
9O+eI//4qPexpEMsQkvyWq3WR4JAnppne5b8C3n03WlUcjV3ZS3Gf2biv+H8/Gge9MiMKUOgBudL
uwUGdNVn8NcJnFupsrGZDotJzDkFIi+fS/X+P0UM6GBJj1sFLnH3NltxB+XIApryPxLLTPzAXgR+
lme7AR01JdOnL324FbavNkqFz+YdE9wBS4eBnnsAsqClVCIJZ+b0Nrx3NnxcbUn7WDJkNIP6PEAD
UAe5EBJxYBogHpp2I66ZNjQnfGfrD2c+C49GxupPs5UxZdxfpdalXppWUTyJwEzIsACeyTnxqhT4
waSRd1+DLXMK5lQP8jZ93uK//Ey8PQrxyiH8V0VKGYzenBe3IM08xqvy9QGxf23jUwsJK9V1ynYD
T64ClG6FbOMIssFpFdZrsBz6zyjS1dkvrSbs285RGFSYaKi2jcZE0aIce3b9oQ5GDndDMXLFgjTR
b5VbIz2lcdHm+IoH9YAScefdR5XePmFWHVlqwG0ZVEAUBQltJROz1b0txr7oelfVbKuKR7s+mTiu
WpVDoTFLu5ZHYSSB0n5Wen6dSqio9/KhT2LiCewYcSYAbyzeGMY7FfncPB3T7GNBwzDmUCfPsLFH
iL5XlYuU6ZpMolaaltWCvnxl7UK802D/gojfatDBniqS5Dm0yf9sBeCghFx5Bq0jq03yJnTvTyOU
dowPPAFIPsZKIQqyL2X0CwR+fn6FrW3GxE3w8GWn/NRboQgJd9290gXjGAcF2/IqcPgsBZN+NUca
JKrI1v3yBog4uEF1GupjfoVfz0Fj1pfHPT+x9RR25r04ynb/jBj7pV/xftqLKsnR9O21ZUlZOVLj
oXdOSJlp89sr7hhGstFMMEe4ymnSsdTW7Ai15fhV6E+JY66Y4ZkBaUGpOkzfNKSMG6+E1gd2ga14
WhyjkyGL6C4Ear77vzZNsvXWGJuja3NqPB3ykRM5AhW8bFWMrWqesF09ze7TH6yyT2qwGmOkyUrl
kEIjbDKfDMQuNcvfKvUWCNYt8jMO/THONIpRgJ/9taQCY3G1quXNEMYtA7vLThZuzo77m3A60JrR
xRIvZ1kDzPqeN9/Qf6T1t3gQGFVCuF+d4e6x9uPbGsOTqrrcvzpomCsAxC01QikzRicWL4TYIVx7
2G2w11Blifgpgn2y7fxAAiMucWNm9STKxjroinmMYTGzlRRxpWW60BaiKyg5C5Q1MlIgNQeY/Lje
TpDhk0clZ0V/dg8SATfR1IbnE17RZdIq8bIYue31QXyaPLf1b4mSOqftAgC+Ko/iYLe9JUyWTzyn
Br5Q5+xQXNMf6om9YZbRZBx/4XOMJbRUW3oo7zvB05NA+TB3QtT+MvfqJACuTPWMjctXVDwZBGSa
59VdL4bpJR2GA+ErX6zh5tmnNG6+D44zzeB5HONTUX3RrlESBjZGefqUiNHEQWjIXYbL5prq2JH3
dEbRhj6+WPLhNvkWKzYcUzjgZZgea0FrpFGSlYdkJt4M1k9Q3sL34PzvIfjBvR9e2OAjbzal9LAl
S7f2sh1oE56dSqOQ1JuREhr5PyGg+p76bdoJqp+9Tx4K8mn6pB2QC5bBuCFiy2jtLWNupeJ9eGeP
srPR/EpCSYuKSCYmwvtPKypY8S/7ccroIrKymbSG+rUQPCkvndsSHhYtBpfs/8Gq3UiTM7ESOKS6
xkVDUzOTO/I/bWB9yzcuVHc7eoUDrCYi5rKhrEl9xluK4ucTs0otToBYURZkNGk7iWZ617dqxTJi
xWE/mp6nzp4+jz58EftU2NWiJZqfvBB6N7D9RC+M/Tc0Hbw5LTnjZCc4c9BkKn0CdUv9fQU+hctz
QkV4U5wTIJs7p3AFLf4bainJjyrDcc9Kzv9n5oF+PHChs0CMsvbkIAf+dAAQeYOSco80AmxOQGCQ
lxb/9EgAzyXHIUWCqiQtMlJFCmZjwPMgrwy9w/oMgs5Yiycd7BeE/0+L0nE2hZ6BXJrh70XJ37+Z
cMw58R4IX7Ck2lpbXCiBgyFXUOsc1BYWLmCd5gTIUS4ihRHiZk03RJUzzTQx0KQzO6NEu418IIUh
34ylTnWuxnICUKPfbaw5Kw1veyTfY66Tv+Fpxlzx+VM1sDRSNi5O+0ta9ESm6zbZmKvT6z8uLJV1
lVE3DvWjST4VT7/qITVHOxdPlexBmbZxEmGzVtwnhPJoFIVojbrLa7eMsZQJeDJM+/wngYoncysl
pIspY9rWamRMR7wOCRKvrglGkgHRFW2orBguUVDDTMYr6sfHyd1s1u9m/ZMH4bPPfO7dSpoxwZ9s
KMiL0th+p8pSWiF3MX5SzDMhKiWNjWmU+pf9TMlJnIDl37KSrDVandpEx69snpGyC4dQxTItUQ6N
wLKQiT7Bo/nzV8dwtH0n2ulSkigJ4nkRS/IrOhd0DwmBfkFykUtWR94ph3vH46X89rZ/RwzDHwcQ
MElwWhuoODZCzH9wqoyObFNPWHoQ35GN+ZHFWPpk6peqr2UN8cmfrRqEgqwrDBp73gVinTCUgd6x
Nch2zHcyCXzbb62/GUhIudxObf5mLC77OHlFhL+IavdrOEP0IYSQqGzYEJOS33EmNX0UPGiHcvme
iVIgV1XmZNGCX/5VgMZSA3c23Jb0vKVzRGtb1RFVILzZf7Qlgl3FDEzrw0GO0PdnqICwOtdhUKO7
wWolnCkC7Jzs7f6CJED++uFMaB9XpmUOMvICdTMnZL8GlqZ4va488eIesc2roemLvAzgQkSLeyae
xNDbRhjT6HS1uqQUpPTByjYXkPSuUVQnp7s3UF2s5/wAOZsy2PMdB20ECt9ZYgGwWaZme+j3mOK3
Gvbkj6qK9VSAQCu1/HzJOu9bcuP6ucotLTTUwyXJx+sqhzPsL6e38EoFTostbSx4QkALh2uwUkyw
SGMx7nB0/odLTRiP3JngYFPvUu1DR2rXv3iy1ITktP2K1ZOppLAoV+dLWFJy6oxZpWeGdCc9OolY
tHXVztA4XOE0h4gl7aTkOhpJrNxG1yxEnXTUldzFHpK/NfRspqYzpp0hEA868sITy77iHJnmNfDI
PlYKYiZfEWf0CtHlgVnOsn637mJkPhcm8WOUpSb95REORbzjcGvPeXKlHtDksBvToG8p0f8gAnJe
bVzUn5lh5+Q/XmukPUh/jVE/bjMtszq8Sr75GJ9R4zHTCS2znv9Rdgy6l3VmwWdMh2KWS3MNHJ3F
0bXlf/knfzPNJx9yVyTN7T4RR1kqq7E5BLNsa1XQ0H0SEWiUVQbjXA7y9ykIy79OcJWhIzTy8Sd7
P27mCE9DTn6J2+ZWCV/Kx1V49AnWxSOOUo9UqeG7jIllluLo9zFIVl3zjkLVoFu63dPKMASWVfVR
ucCiMNFqV1tEv28DXjVkhTKF9Gxgtys1QxjslVjLkONlTl3PFOBa3p3cesL6rdE4yRh04ENunLzL
ul0558jbXMMmElBCg/ac4AOlvl9PCjt+NJLGh03fMW/7Odg9Qs7jv8A/28yRvMgBKuiX2YSf4QUT
P/xX7dVuavUQZLB1uLc50FOPsAxchFZxwVyPz08My5KYQB2W3MKlkS4+AXfKr6TnXQOLrF8uK+Yv
IZZw1JWoKVH7V+fWtE6Va7XI4yXv6DgxmHOxUUg3kQ+yWnyBmEDE1VPC3SxgGiT4+KxPlsIK4UDs
dvr+8ZY6PkDe7Ei7VKRbXJT1Cx8eHErfOfpZTFlMoH1AethizViImAkyGPbKpNgDjYHCM0QrehEp
yFSaJT/CpXvpjZFS3suCWw26ltdCJGMA52RDwAsGFsFqaPcFKlYorq2+h3kUrhghe4mbYIEohqSq
+SE8TxbdSul/l8NFhkRyeMzgCjncBDTQBsy2WOJbMZFlaBxH6uqL7pIg4ci8r7WXvTzljFsOXpQB
kCGSX8p0YO2OLP77OJD2W3VssajDS+B+BXS1G//4eqFQk6e/D7yt9an5s23dfw7cZvSzGWaxgyP1
d+11OJbq01Wt0kNMEmOr0Q7HkLxiO6a0kJjcTA6X+r1dCKmJ2Aw2s/EkzXD3zrk0Rt6rSLYHwByQ
oN6aeMN5nCUJ4Qeziw+2Oz2GSZ19wCL7fPIQ/874E5jETG0CmtI5qxo7JIsAp52ZczgeEo0iLzFm
vpghzBentU+d8e4+j4NGA82wH8o4kiPnjitdA9Dbk97+TfR9vHbrdcC7PCbX5USaNC3hkxAaDASc
RMEHBw+A+butqQVVg4LtPWSgGKF7ueLGktU5TXUtUQYRSnQxv9f3y1PcKFAm5FKni/QYAEP9U876
1PdcxS8Ee4F1G/anmLi1/ioMZcX0plb+zEliIUcpdy/phdjk04ZDJspzbkBU2pM/nWhp+ZKl8ul9
Hbt5nppUzOYiTeGInmw/mxX0Ka6OFIbKr3pkPKsvGhZ2z6/sNhLD+gx7wiqyedmhcUJJuzFQtwqY
jN6AJizjdT5TvIBexmQ2gJ4Iidszm0XdZS7UzmUXyO3PC6bo0BoM5puMO/1SOCQd1lZXo08OTPKz
cjpxrqEmvhWvPoaN46iB6XHvj85G7VuMp0ZrqLcpz3pbGzY5FY+OVKuNhHcdgODD2264LbJyxctB
qmDANZQsTEa/xTxOwzfBhB5Ru6e58kEGpPQBaq5mto1qiybzDCJJenR6ruYws/fYoNUJNy8GbsSp
Ju2usS0vgUJlPZwlsvmkhpekPGOUysZx390xAk9p9DuBexo5HTiAgE8+yvEY06WCsC4Bmh9xcF01
63qcrSU9aAMySpXevJLMmrtFwxsauEf8BvqTrpjVBf8Xr93Dy/EDgltfs2OPXJitnwWMSof4QJXe
aaidSxQf6wzxLtzywSSXDxIRDtDcTyHTkdKXVj0VV2ofAV+fFUGh9a7fJSMy3ChutA/hPQVbJpzI
ZJGs+qg00QBbeH/4whBz7DZYzVhBGXq1VJZKgZrZ5rhpsOxE07s4pZZ94UQE4dLKYwBDKJ7dJIbZ
+rKKloHOvrrzr7fMVSGODelCplbWApWWnGmXBWzIKqCRV8NlJLXhhd7WgKb0PTbfkVhDelMVoov2
QTFzRfXyFkOlFUM5IahDvuIzyPhVBJW+GaBVba8JZNPwn7CaxP0PNy/0jIOYljXQujO3O+l+HOC8
Xk5/fZiAvCzi7B/146Zv9myAGSwwVR4sN2Cg3fzgRwhBqdXLXmbSgpIuAifhEDNdIMy9cAmCeYV8
qEgUOTkRSlXWH5hbhJPU8qziCXIBdVW1ZXA+uP+9Cw+pSzkdXo8qqBh1EAUvz7KQm+VjOFwQpjlK
YhDFXW/s8pP+eneojbxmofPqFxidv1ps8fGCidynCIpqFvMKI657vUp8pD0joVpI0yMlKqQ6lI1q
goFUtcL9fqbzancnX9+v+2gZarKTh24Qt0aGy9rOqe88BFIRHK4hjbeYCZ/wnihdzXseWJMk0uVY
qwo1G02Kv6r32YjT63gP84NPZLT5/9hXjT3xdfF6ld5Bg9U3/znh9OzXLToa+1jdJDXC9zK5jLqI
lVGwL+MstHpk8lxpQJOG8WI7y0mX/pSATHK9PeL8lP1Lu2shLpH7JmlqWtPdTmZ+axI5tGn1vc2p
51H6cq+2pNE+MV1eiFN7Ar5NXAgk9xp2WG029Ohd43uzUdEtGwSs4GyEkUnqik4EbRJoyUVg3h15
keNI3an05X5X2eEHqNiWnzL3cBPHJRk9E7IUuA4bSPiiL1aCDypij8SV2wY6ItB4gkd46qPMC0ke
zZIoZfDsql8aerHhSMorAPDHF1MWCYT/UoofPFymY5c6UttGMUEeXCo/ClvRg3XNEMBmETLCHKG5
6cjF4YYHhEj6PllW9G1bDmSmXgq9afVKcGfd4Z/wCM1FAxOeaDgNca+9UQ+ByyEQZYwbdNDaRmqm
n9KZPSX0De0pB9DzF8oLAyfuRafL2sRMAoz3YZUkog5puPym2TaV5iAUDLC+B/Ybvu3XoqDYCnKU
jvRSlqmsLeGwAeGE1XIGvinrUvN7FNH4Qwunfo+QDg+7eknYL2K2NF3a6cclkrxDZkwhe5Dui1lo
e860QpDlKfxUeU6ygrmcg2tdsCUpNGegbQFQXy/U7MzBx2hxt9IdOWed7eRIi7EgqN6xKYiXSlXp
s2vDvRY0YeSqi7c/2Gl/OnkJpgbtErUK0d6mKn2RJDS0DNaxR9NztbgYOoJ03czbfgtVxBJ1/pXR
dr18IhKTnnxHGThQkUDEocrkrdZegEqKRPLrmkcTkAOW5CUfrM+lhl+OuuN/fRc7KpmEURWZ4/f8
2MSuo23spaCo0gXXVWRoZbrBM42avOj6mpbfoCK1adSMy5DPtAO34n0EPckTtf9ZuakqgnpffLKD
1PuwQn4EANgol3HHWIAgpNy0+lfmwlSBY+8l1fQix2lYMmJvQRFnc8CdzRasHo3R3aTtfjvPk/3u
GS9qL3vzW8W8+VjBd14tSijR6cMwBnAnywQXo0HQg19RhUKmrRPwG8t4fs5gMO6OOX2DLUHpOZXS
YLarQ20VhrTLjT/fnTOYuARQTEWk6TaPWH0vpeqn59TcQNDyxp35PrcRpPrV+UEoXgLan6ThAeXY
wnvqqROnDc/uryMYcg5W0pPz5Tu7o/C1koprTRkYxB2Yd4dyv6wOdK/paVS02g6hyfSRMhNtIWMO
BUB+h/vdxhZlH7d5LcJfD3DzBIuVBwzA4Y0ksHGsKm+Lt35GDA6IL14/fnCSvuWqtlg6sN4lVkCj
m9lmEA+iKie466dneHuDbv4NJvnFvLyJj6gQHZ7weHjdWCe3RY5qYdwA2qdHREYduVUYkFxuLNQk
Q5Aiil6p9E9vrwA02sOB2INpBBpZe1+4hlu9ocmT0nRtDJGa36c1WMvjIHPMx7zHfWEOaFSXWun7
zz9/9GeyMJ3yqIz+EGynonhZBaBRcELtSvb6JXmO9Aa+XPS6rG9w0J+BQJChZsmA1ouOsBbvrnoB
aPNJfW2QbUjsKsn0+GWi7Kr4Rj/ngNjaHlUuHiDFz8jQj3z1RVSCXhLAR2hObBVCLCc15WqLMM4Q
Y28X6HQ/83chqtO1h35DhlrNxHNM8GEKC+I0l7rFHSl5XbiyFXXDvxqbA7TakC6uddch/Q5fgbOb
EHH5IPvyrJCy94VheGqc60K7T3EUpz7KniRochQiIP5ynFzmUYX8lR/DU4jQzokyfvW4GDxAyLuN
E0v9ZhOEiPD+TRgWeUSyzYYSHuQMa0WeJiOumtixlfUlubVZw6xA6E3lnPPs21h/GddZb70Ox+SZ
8n6zPHTPFMhSFoHnqWLGBv9mZMSyUTv9Sc4HRP1tnQwIwdTUt/ZImTzlIRCbq+bsY2F2sxMw1rQb
2KYjHLrVhFd74zgfShYBVBjcCN18ZBHUxheb3dY7Zt6KYKU6ampv59nzUsMHWSWJOgueXyQdVWaL
i7Zu/IZ957ruDB2TgiJz6FOaJtDTajjlYIv+DsgOmAIoEukeKCWAM3QPVDQ9L4My/ypDR5ZCNSyO
YCNJuHAIniCM8X648KX1/8/1MobMiWAjAUh5ZIs99i9J1I+vurQjrK51NS1hF/7V1STU9bY2Seec
pXYQXoNUgyKmLVFyNyTk5CDGmjAvv/1yptMHqdNr/ypWSM9nMahHR6gRsnPYFO7CyzKKZvOJHo3J
6P2ORNV9TfXUqaSwW2CAAEZpnFzLOIFWVsMNn1NdC3sn4QKEVHyZ5f7aD97cAnpsFn+qjhzPeHb5
cYdCcBCsYsXOcaOflZT4x3WnKU1L+Sbe8PZY/GfiP6neOOPy8FTGPIZINU6zXknWs9Yvz/2Af679
+VF5fMvpQkkrF5FCPzmhwnJKjH0Pf7uGIG2DDGqOoPmvbY+raLVVlJXD+nn3hACCG52rtoR1VgE/
a4xafAMLDrf+71ohIc5W4VaPoHZsG8pmqbIsHRtElkfB9K8C8TN2MuHKXYvxEoSgKnTEMusagYst
Ex04pVUOOFQh+eK8Vx9+Z7lHEo8j+sIVFPLSEE+haRWFlL3xU26olq6mpEPPl6JtlHQHmpGfYd5O
GEc6C2Sh13656hvDDYL3gOkkJmJ3bwelX9dpuikNds4BOsjuyiuCWLrvaSeS4vNpH2eWmKs5QEe8
cO1gBsU+Jsdk2tMKAFNUPyGSu/UG6CDl33QzPn8GOE0md3BvU43rTNTQHWFBPfHWvNR3PbCPDyDH
clbl04zex5ikgMWiZxJY7mCoirECsDgxeaLzcT/uIubQNYA6KB1VlNtLgJ40kPo6eCtEA54MGGgE
ktU+4ZCcwYhHFEAI0k1nP/ET2c4oyjbovNKzTfZyxMtJqL88cjTHO70HtaSHWuSoRhZTSqs3Nq/L
NNTHuLtOcmthZG3N9oYfXWu6gSUpaLqVO6FOsX8zHXBROsTVEysLHTA9Dm9FIMh5YEKHzctmp/Ji
FQQMpb0dOGTMRPs3B8jqTE7IIgJ3qLtVf61NeD48XsuvHXpd8/IilywbNbUU/vBo8uepnc+CUa98
+vpOaHbZbDPIqQLt5poHeE2booNW5hlQPAP38GrSVHsRvlBvyCdWuBFzMBG+DYCRsnBF2bo/pt87
hXGFkKASgnP3aav8uczibmUOKT99yw+Fg89dPkusNNGyDDdFcJnHrl2U/dalhnbYK+5fFtki0VY1
Tp74+x8TlI/HrfQ6mO/V3c2ghS7eNNH1y4QgX/cCGYxkDmg9p2yNARSYgcW48rU7YZvzjqntsXR4
FM52nis+WBiAMm0wSo4YH1AzFiDKOzLRbtpwpyFtoFbOOx+lv2CJU49PKWtC7A8HtjgiD08kJmi8
ViwmzIlMGLHzGNRBjj2DDX9uuwJhg9zNaN76TTOQlNLBd1+aP+FqjBa1XffqZ1/pSskXCASvbsBg
pM5kj7MO1QIzOU0J8mvR2GovZOqgQjM79RSbkLqObkxa5EY87JbDQ62aGK6AYg2HnXUInboV1Ed/
YrstULMLAFzzB8gchQaoyt96amVPfDxg+11YwgTtOr/UySUoEs24L8NMsxOSA7AuK4+sv5FTy7hZ
A/AXZoQEyRcy/W1PS2jrDnptvWqWvdcSXbXemgIAhnjkMJk3oYzqZFTvpoHj6FQhxzcrYt5CPgdj
GpTrkNq18IyFJTjVqF8I6UIx5kCFgGijbUZTe2uBOINRnvFexOZw/Qg0h1ZtwP05PzCa/Vi1eT+j
WrOJ3CLPBP4iL++2e8iQPBPt5VQrv0OkOVfdnqycYqUy4qSfc0dARF50bmuWROuN9xiNyKc5Qr9O
sDWIFp5afM/lbwIFeB9W+WQkH5QJnLyipj7QTMX3mn8SDqcMqaMiOTphQ7Yh5XOq7sSPTECVkeuh
HVlt1IaP90HRm8ME2yiNJjhufpHVh5kBz/BffD14CMCdUZBU+VdiB7gc3oOH7/Ugr3a3QquvaCDM
rwuhlbpsue2H0FNpVr8tjpw5sovgI98Zi5ci4NP4NflV5CsGIoF6pEU2qXWfN8a46nI95UeWWbn4
Ii39AMcuh8wNLpesml3MNufY8OjdB5fK4f7lWMXpqO165bQhGOPQZnCG6VkGsQcG84V7AhsVmP5w
ZzHNI9obPRU5QPlTSP4TYiUrFMTDJDDd5O0iDRA5oPJ4gjWOPsJ1bcJ/cO1p2wUUzvVd2R2Q+JmF
MFLIE8OpMKchBnkWWgf+2mtlJL6w365Dy417h+xvxMINpFXcACj05LsEA0Z2m4RqTe4koOI7oLey
6iKQfNievhr402rId7MblLqyn3j7HQ+9aWVA40uVCHPQ2qGAg/cSi/ZwSOFjcGRiDzEj13R0G6hB
VXTNlg67RaJ27OaDIJk8vQFLolwT6ABmPgkUS6YqGdnycu5ANHEUcY3UyH9SmFe0MgEcPiKLR7LX
rldJyASyfo5cJBpnnowywsEcYaU4WyczxtXj8k99AitDphHMKDlUTFQhL9lmEtbxJaYvTIvK3Kie
regQOTccrSBLeDK+lYzuBYw22nQnIn2ZD9CCA58Cdp7QrVNeFnuGD2rDOGyeuc2arKiX7MACq7YI
hi6TdH6avMcv4+7Mgw4OoaORkP52CWVAXn1jiO3pBA9UZknvh3o+CdF1AWT1Wgl2mnCiXv8g586N
VxyyLApJZBd4nVBK4TG4OQ0qc/8rd8oU+RIohZ9WYWxM37z+ykFvClFHZi+OhSDdndEDmwEeDYxT
Au17SLiIuA5fn3nbXBq18zVhLCka6hB31tOyOhe8OyAVhlDZmvx9tieFY2CJTXwfjN5miaNpHVuT
3PaWQ+Z0rPP6HGXHYqDhqG6s6Ts8ttyiJhrO/gZO3mFF679BTC0J65DyFMIR+1jqAKfMdRBdZUTi
0x60eGhK6iIeVuQPl6kHSPbz1WZYEcEPTga0pN1bNrRiA/lQQdsC3keaENJczXn8mAXpmK1llmGA
fa17Mm5LpQMpQSNi9+9LxDouHA5OBovJQ90WIQuZQ4R4QuBdXwttbonCVG70UA16ALdVYzJncK4J
BS3FWEFdpacbO7i4EWlvjcDL9eyMwKGNNQ0bTmYgcy96PH9YyZXhTbEnZajLELwORsrGoVxBjpwK
V/6xHRsb1M4NtJfutQhHK2v7ktdtZnc41qfRipKLEAHSEFMUNz9JjjI/K/3wDCQGcTFfvbd94kyR
wZEBTXutUSCWfHa1L+w+tCOFlZy1py2aBOS+51wMBkvHmrpg2VpVScaVIA9gYXofZu7ULpwBiNO0
6BL4k2X4DCprbfKtrMnPWbFSsMcc+woDjKqOsBfniKw8eNmNlkgc3JDE8DvGK5CHh37LIkbRHa4P
etAyP7tUi64MVBRokHJ/yJOFn/3HBnMUuQ42uABKn9rocMWCkq4EGLP6eU6x9M6QGivUeeHtY9oW
GcrkOHsjieAnIJU0OdlLWGJMhixDkefdrRk3axXI8Zt0RtDuL/W9KbpiFRoW9AQpARfLk7KFNbGi
rGQy73TRQm6ciI2EY9NaC6KunLMj4Pvh+RNGdNlHdwFOEsPBnnwRsfdKFkFIJn/cJtuIpQ5WvSQ9
I3wWtn0Byzcck021jdUPc3TpHvfI/lvaeQRYV3cwsV7aySHqY9nVCJ7CwuEMUZ3VFnaPq5/etrPp
/WS1SlgCVm/dvlD6nmame5VmNJtfdmExhJGkGuE75yPIKR6JHPVW+yYbhothSA8p42Xbj+BJwxtw
HGrJCgbilpbFqOVdlSFuVjqaB8uvwCcOq0x4Nc1j95C4BjzOkgrp2jLtvkDlX8VfYRpSReGvoLUO
0AsZA2zuIL9ocH0nfwMCsMHr0CUbvfzJ1RqfyINFMeNNKG/uEbsI0LixIt2PoQrv883VY+19WvO1
a6Mg56+jB+siYrDFztFLderF+Wlxl2Zo4QeO3cg/Nn300m0iyU1tsCAbnFEhUIDt/NBa95nh3VyN
oS5FBRqFxNqYOhaSeSJLa0VvCI0pl81E6qfWWfuMW9LnY+1ZnMVsDqpzU2NAs2k6HzS10xhFnj+w
Lrfy9nriFrvoN47hEEzbZeaezYJO583iNL5wbdU41XJjqmOihZMOQc1GgwO2jLkgDDlPZXHPUkj4
pcmtHTVBfdjB+bNjKg/TrBWEALtGKJCg9CdAMeFYRYdoQTiyxBN6TuRbaSNkbxiYUCNfbw0w+Cak
phnqMHUoeNihXK0s38EPgdwRMeNAIqYhqWVWeW13CKNVAL38UyZbUY1wNLDmR8K6rP9oS8boX2NA
b0eOOpt0UUlL9oykB7Q6mlydJl2ZxvIyNEzhC8by1cH9Jje/w0RXt84Nc9MZhpwuofvGV7hVzcrs
B8mxzItr4aJOCF0nA/utEILVv0r47x0qDid2cMKKfWCt6Is/rTbtAWlQyV7PRIlKlBL44jSA/zCu
mqvIpve6+dQ4GdNEtM/KrxHnod16UKWbjMPidgIgd73RVsO9f3S4wtsG0vYLz839nv0QJhUpl0Km
DLG0+kLjvyHV6vlrXrn0bKirHJPazWfDvI46kJhWG/mLam0uNkZYdtgb+wEQS5tsGoB5re1ByXkn
xb85W86KuGw2Z2j/b4MNm2oyRs4RW4jmT5X+C9a/LKn9h3EZFBi6B3j410VxkslfjsAdB8mI8NNt
t0mhR3kCecflopq0bwUpRWLhyYkAo5xI4znLItINgOkQzPDj18xZkhMUoD9jLZR+AutJvXmU0DHD
52kH09sZEiJ5FP/9ZGY9uOJTHqpOILOL1fFJe68+P3B2PYK+wbZLVDSzK1x7H5anhFl71WXfa9E+
Lt+g3w9opm7KnpxpJ8U/kF+RJ176JQrFrxuGV/2Oi0uWIC1vPp5VbEHBE6Mtu9o7anbtFRNjD+oH
KsIjg+vwH9pNz9MeunLWYEs8/kBKUG67Cn0uiGn2XWI92GCvG6GVH41Azj0YhCovCbVzUuIeZMfE
D1kAV4P8BfukdeasPUHCn8rYVLb2VYpq/kA0K8Z36DreRKKqCQESY+EU7TSMsnSFy0qjwC221vO5
dDvEZsJQXGzH4t9xvuTXdL6OEkJUjrlicX6pGVNGjDDvaadQYrp+Pg7V2uvq5JyxlHbek9y0UOAC
FvmdPszKFvAmMumrlxPkgskKt/ueyBufvrHlMrJmAIPP3r5DvERObTrb5c81RQ+I3o2IuSNzXCqe
7huZkRl8vTBpxPvXF8tJEVgFBIafls2qCq/tid+CHeYsqBTw2RI3DuDZI3zAbrmMZa+sdBtTGXrn
kLSoRxlu/SrkFsGgaA+lJXbuyrS92UIH7H3KJraPhPEMQfbtGFVLtLZC1AAmwP3HtZ8blbLjmELK
3CxqnsjMKINa1S6p7t9SXYze5j2v8JH6Qz38++dbmIKStioY+d78xyu6nvrOKJmj9uEHViiOHFRh
iV3AzEXEmyKCcX/R/SQiYldfFmzKo9STHQlrcTHZA7Av1j1IvYj5pYhbS77Xbs+zP6lPH4qmT5RR
7jZdiwnSxBvTb27iskQvjwmIXaKxq20mC7Sm65OW8SItPkNwzNelS5jZrVtiuFn1+JrZ4e3TJlgl
2zbi2+aMD6F+4J5cxZZe+YIILjzpyfLaB3TYXCecghYPJlS0Nl1CkBy2+MWOWhBhiLUKGv4IwmuH
DSgoLSU1Acwao2NrYij90OtyYiuwIUO6II30Zw+a5Vj/JiwTbw7coE1MzNaZA5g022GO4R71HsoQ
Whpr+8cJPFa77ftMeOUfkaBGTdWY+YSCuLc1ypmUiAxS4WOkZSUuob3bS2mTk43LOnA3P9L3gZc6
nGjbNcjnk3ov/buBfWQhxnirhFF0r8pAniNH2FPYljflNM0ry8vkxYrMleyIiwL5ZWhvJNv5IzPV
uhMsP3zVraZfTviA2tcfPgpNw40W4xJ34GytPueHFx8L7I9HvKn9HXZy+NtF2kY2WTjX7raBy7hx
OagHTzFhUoKpBtObSiP+ffbWuL4eKufhMBJtLQX7OLXQgdZTAVDyQVOstOM+E+wGNkg/Jjtl48ju
eiJ4Sk6bawTDOEpvVo1hlqqX6Q8VHGCI7YPeI9luSvuFREj+/88ZGor1tGcln4HVj2QeOzjT0US3
GATirlgpCzRXLOKIG2ZvOppa3KK1LiOfJqUwd5ugOueobKeMH/tiCMa08UO6mFUx2RAit/cxBJFa
FEKW8s5sNoRFSf1aVpT4qnByVXikUGa/ijDiNtNuW1VfuIUnx3p8XiIVYQqwuabd4fNlDKHF0S17
4Ftq3lyD1yRJP+KtJM0KiPXjWUfAA79I9Uvnhzu8i2BpKOujj7WCpmXSzfrXimm1yCJ7Ip63HGuh
Z/qoPuXmC2HD7VErMaKoGy2tDXbQJyLcHaIowpN8rAiTcZhsfkNrAd4vnNKxlj6PvIq/MXWx7oO1
vydplsjSNP3UHPOfsK8XxJSV/Avw+rrxL/j710pI4djXP3rr4S+XKcNcbqKjS4uwBdnGJ5poyfxc
WuByvJVtUr5qPb3vpgwtEXiWCyEeet90oLweCXBDmMcCgw3gucnitgdZ1o1OH3ndBgMYRHVCNqTo
hrla1Ao/840RXe6nxhWs93KyVuIzNZFDFjqhmtr69/oRP8J+G6s/CzwyoKY2KEgK3o2iRl+O5Q8T
Cp3Yl8wrEpH9yDk9nHeZZCoYk8/5ogWU8RHhvDa3VUgek/exMPfecNDk1wKqbw8jl+6P6x54Yu5V
UAqLcIBveYnLcHlVUWZ02pZeXdmxp6irgJ+Pxd0IY8ISotAiARZtsZeJwk5kEcQ78hn4+ubI6zTj
Gm5pFCCd43mJdx8fYvBero5d3aEWY6B7B9wjmTmxs21FBqJ91r4KAfr5M02BnOpxvbumVDEb5xiQ
cqy89XN/OUObcXtCpqGOv0on+T/2ELEQUFyD419YRksxGPx1DXS4fZ4StycN6bLyywJgZYJL8/nw
gC1Soekeu+9yaFKpRIomMvMf+gH2HxHmFVFsiGTohkpKseNEhNDi6SxTkQND2TddGYTs9trWM/Ru
MT1dQDpIVRQmiBApMLFr0RIcSIOGNqdX9M7o3lFRHCpPlHl+wQRacaSpt1KB/c/+FzZoGnL5COyA
rKLIhJOYHePuyVQ4d7fNkIiRDLPVCGC/ErtNHHLzgbnLZ8EQnZSG73FQdi8SPZAqBUJED54uo1vm
eQqmG1aVXTdMB4m2idVFFU7yBerZrCw+/LNh7qWDJPxW5pdhP4W5qRgLb4K7lOSXh7wNeqZaO+F4
TKynBgz+Uu8dklrzK2E36ONgRGBEho1Wo48sweMJwaObeNfw7oejWcAKA32kCT3unIknxkkbesnP
JjoJPvYYhmG4eNLZ2cJNYmkb13FEyHa16dP3zCKXGyy8ZhBj3k9WscOI7gGdqfcHLwt0gbR/MXcc
bkHr5TD9ulBQlTj1ssVDJThEgOVKym2zWAOdQtV9ZEIZZ3ebURpe/OT2e+nkoDKowSKATNGyA7E4
NbTy6HiSwUtAS+U4JuysxNHhSnDnqCQKyAyPqypZLheMhsLVxmWSMZsK4l8EkHKs4mpUJa4tAw+5
qnJ4bndCodsWv5uvTj/u93M7Zb5PvvV2F58YvnlNuKlHUjNVPLs/RULnO+SBiRWxA5WzwH0JqLGa
svZ3HHK2/ycEKv3GPcNOABy6MybL57uR6dKWFvt6ots1wmzLtJJyJppOA5BqEZeUHgfRrtfonxaY
1eqhdQgHXyX+F+50CrjZQczHUbzZ6xwy0ZqD39q9vOGuGtb0kXZZ+ab0Eieg4DaCs4EWGPo9Jptk
PAiP7FHfRVR/IM2npN21KX1CrWx4MAOMuskKdclE6vcoyeEdvp5Kc4D/I4ofyluYXFZVAN7MtotU
1ZRMcuzxswGI2dbKFZWJgpWGGmGk9udfy/+qjk0YF4eyJtr1Ru5fx9anDxOSMtlkVuxI+o/p/S52
0LCT6IBfVGe2IDh5TikPCeAGM2M7avK0k/QeHLpx6YbFhLFoRvL0q4SYirrTd8AoDsQC6dLLVvTT
utyGJtDnmdw4b5Yswgf1g//MdOeC0AXaAvoGsMKgmqPxgOLL4vsvTVN3/LZu9gba/P0Y0M3JZ4JX
6XugIeQw33lb3C0lD2fDxixs0YFdSJu7k1KWf2c3Fa06Ae6buUzIEGW1IZy/XtbYTiNgcApu28ma
jhMEu0PQWnLhKYuxl7KfIPK4HEC2a486Bh5ihqDtS0lP59scPT0G2UMweD/1c0Z7QBezy9DJtV5l
ESuCfRm4bMITG1359hXXUBs1UY5FC9h7tJY+kmD6Eb0nQS0eZGafSYENzPPSEJzRBf1w4HZTQOBK
cioKZTma5cbdsqtKb6L4RP2fFT/SqONdSm6LxXrXeCnIPwhd3s5E+r5V20NqgmTr0N4JfM//VAiy
hk2puF9HLHlvLUjFrDg/CNvwPAJmBpbnlI0VJOUUm75oLosxXyyobdLEekwSr4RWqL9ahXzYc/m0
CsAlANEDaww1RkA3JkR6zmoyT0SOglI48CQiAizDFccvCO3qI1tPQgtu6oCsc/SbwOTGpRJ8NmQR
PQRz5seybYW+NcZe3x2TRyfaREof5D6FUD4uZUoHLdLS+vNoxDkyEdGdThLftrJXYabPfJvUjND5
KUt6kdrWdsjF2fcTV46shU3dO+DjHHd1hxRemjzVbPNrOvR5x+FOGcg+Ul8nuJWGoE8si/DOnfj2
t4u0ogfQfFd9cSlhQXW6cr9eD9hvnX1C/0z14kl9GE1nDDYH91v78GYFQvkx5//GFFPPWlWS4q2V
5M5/86zFRefukmIftzs0zP0sNImii3d4Si2VRK/eE9QmY8L6qs+0ipG1ii0uZkYooffpL06sKwhI
N+13IcEJxHYGamBim5iRepbyo2I2QwnEGq1llqKYjpxIflbfsLokLFvA10UKv9l1Ozq9+rKOG1Nn
63xv0+Hs36IDr7wjOUdfqKUppin4HiwGvNMpp1wHesEGU2XBRR6u6Cno7i/37YJtaICP6wCOj3ui
9cI70WfFbNCpQe5diso/3ihwh6Zf+BBH5OJ0aSL7aYmvtEMK+LUJSzkf7u/oA1mw+L2PspTTfxOn
VbRYMvu2+PSLeBMQgCen9v4icILx75qJzGGBoRpBRIHG7hAS3LMDGKxsmmXw3MlbyFjJh6KOY3Zx
weTS109eGyxluuaqm6J7PkzJ6ad712Dz+39hQMu8O7dmT7duSE4KB+v+XB+HyZxqNWZBm6EdvHJo
uo+K90WiyJzJ+bbOSKDk04RGqVPi029oy9lslOxbF+XBIzANz9aP4gl+hpp1CTOKgIqg8o0nHPMg
E6t/EfKKyhRpCxQhOJtZh0G9bChcyChvohROmdr9agSoFAMYtfpWawlqiynx8A4TGi2JzsFn8hXq
vNsPOCG1vJLHWEXEw/Z9TpI/lL7dc4RlMIvDVFstOvGutEhPKgOAatuLS4ulqsFDXZMfJwH4Otqb
3AqS1RTlowxmFTDw6xbFrt+KGm14SubElurau+Z8bkmaVrTbvB3x8sGXSjYmLWDW2JbsMb6ktbvt
I5WJZW4dyNiOJsswdENjpRMuu5H+2LE5tHrIgHkZK5As8fzmxioVNh2sGmutH7flNL2x5zAGJbyV
NXUQwmP/7C8P+wvZPEu7GjfRbS5PLmmZt+3Y0Eo+CWij/fGwhQXvbEb0Bk82S+YOW5uCy/HlNnh0
lZOXvnfsn1hZwRFacLcsD9FkfzkcqR2JTw0myFZuNKU6iAKp15S9QQAgfKhfmCcpWRafGE+C+HgR
NgZJMi81lqV02+uMJLnIcmHnZAuf9ZojZeG7tHOMbKa4pqXjBAm8zkJvTXbgLpEip1mhKl3lb+Ds
uucvk9aL1trH05/+U4VtzT4w8h5+Sqoj4dAVRj0Jm9vtHoc7+9YfukKpxK5G91oHH+4w1rLMI3RM
gOfohwTIW/Ig4qnjVSlsRs5immxlAC1+VT275vOrn0AIHsGymUPsuuE6QdYAPDN3aq1u7svNWijO
oo47GLGPEyhr1/rgfjmvFJeTKmgrpzsxICHg0eVaJoOkWGj2uJeDLhvv1SJUeOTnP7NW6uW9c0rb
Fj01rg4dbA9MiJeAw9sHJhQ9he3QaLIkWP+3pI8eySuANrR8TvO9g3PiSgAPT8mIO8OeEdybsl1H
EVMVSo75cbcbSz7tXFwFrUt0W1kMpbwvLDhdj8CDosXSuAQsQJPLCRxDEhkSuHym+r4bGYLXBFMs
xyeOVMnr+t45czpDEcSRsMCDk3xT9sQ1jgcj4lxfbHSU3F8gJdXih06TX/nYIKs0L+n6VRFWhYd1
zGExpz8/1s+WvaioRaD+ZTZ6ZTwEV92UHYtjXsEchAfwarkZ7FwaCeCUnO5iz2pwly4itTkutrDh
2dm7LrofAAgMRldIDXcKBdU/O+SP8Oz15J85Mkee/cL6j5A1iwUyEFLuQdDfBbeYLXz2cBOvm3WF
esRvh37ztXwp/OvTwhf83moj1zqr+RU4jZO1O2hOt7lDcUf/dYCoQeHEEFeNewX5aecl8ZBISZ4y
56F9uITekHV+FqLsASbDevTMRRQ86kMiSLirzDj138n2vecTWU//EVzM9Pbv+A6yhA5XWQjsTwBm
fqeitX2L/skCwSZo+zv1hhpG9A0fN8dsyD73zYv3Qu54VhcpPBZ2FeP7aW/cNUOYOYsUMVMfiOaA
hs8W0rsFbcC5Gg7r5WxWr8KnMnBu/zjua+rB/FdQz98f8Ji0oP16myW1GWRcgC4abM0G/ua9lr4y
ucmiDoBroadJPBbgYQhgtoqLyUgeye3Y42joTuBeOAkKLysV9CnQCuGsFFZjLZiKLhV1jGFYMKnf
VitosGXZfruUExPZjOJvQZArvWNLJz1Dvebn/y4hbjU65eJJV/T/TI9bMwYcZXp2iA9x4uSG6ize
FdPBWJpmOCRksR+xMeUJDzhEVTm1zNhsUcdeGk+lg/gs2wCY32zeyTu3YXQ+kj8YBRjnzoU2lWCF
mXvbBzcrEasmzy37648Ahwpla/qiDVvkOacJoQEvzhAR2wu8WHbPvUfIvvMcZVV/ede4e4+UF78D
oh+8aWr2wiiI2jIowcgVz9/6wYJAzrxGBwiIzwHeYWbILepG1+0JxJJvYWNcaxgJDsKA04TL3OCT
kNr2BpfXHLwYLJw+WW9++dhCQ/w9Scym3GR3vnPVMlvCMQCa8ugoOVDAB8LrDgEXPvIhQOz3VnC0
IiI4Jo4S2XxfFdDrgkaLxKqdTQSZpbiyxkogxiUC/DW1+n9BQeKBp21Gtw3KEOCzz6K4txwZmAaH
YfWZq2eR6apxr+q5ZsBPbR+PFyzj/509Ng0HZIvWm1yR36m0AJfCXiEb0A3Y5c/Rf6Yx4eY3xxaw
r1b81aBZ
`pragma protect end_protected

